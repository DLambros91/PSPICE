**************************************************
*	Name: Demetrios Lambropoulos				 *
*		  David Lambropoulos					 *
*												 *
*	Date: Sunday, March 1, 2014 			     *
*												 *
*	Labratory Experiment 2						 *
**************************************************

* Model for TIP31 BJT
.MODEL TIP31	   NPN( Is=2.447p Xti=3 Eg=1.11 Vaf=100 Bf=208.2 Ise=70.69p 
+ Ne=1.565 Ikf=.9743 Nk=.6134 Xtb=1.5 Br=12.59 Isc=11.68n Nc=1.835 Ikr=3.86 
+ Rc=.4685 Cjc=142p Mjc=.4353 Vjc=.75 Fc=.5 Cje=188.5p Mje=.4878 Vje=.75 
+ Tr=194.2n Tf=19.85n Itf=164.1 Xtf=5.945 Vtf=10 Rb=.1


* command 	collector 	base	emitter		model
	QN			3		 2			0		 TIP31
	
* Resistors
RB1	1	2	2K
RC1	3	4	470

* Voltage Sources
*	+node	-node	model	value
VIN	  1 	  0		  DC	  0V
VCC	  4	      0	      DC      5V

.DC VIN 0V 5V 0.2

.PRINT DC V(1) V(3)

.PROBE

.END
