**************************************************
*	Name: Demetrios Lambropoulos				 *
*		  David Lambropoulos					 *
*												 *
*	Date: Sunday, March 1, 2014 			     *
*												 *
*	Labratory Experiment 2						 *
**************************************************

*		Model for 2N3904 NPN BJT (from Eval library in Pspice)
.model Q2N3904	NPN(Is=6.734f Xti=3 Eg=1.11 Vaf=74.03 Bf=416.4 Ne=1.259
+		Ise=6.734f Ikf=66.78m Xtb=1.5 Br=.7371 Nc=2 Isc=0 Ikr=0 Rc=1
+		Cjc=3.638p Mjc=.3085 Vjc=.75 Fc=.5 Cje=4.493p Mje=.2593 Vje=.75
+		Tr=239.5n Tf=301.2p Itf=.4 Vtf=4 Xtf=2 Rb=10)

* command 	collector 	base	emitter		model
QN             3		 2			0		Q2N3904
	
* Resistors
RB1	1	2	2K
RC1	3	4	470

* Voltage Sources
*	+node	-node	model	value
VIN	  1 	  0		  DC	  0V
VCC	  4	      0	      DC      5V

.DC VIN 0V 5V 0.2

.PRINT DC V(1) V(3)

.PROBE

.END
